��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��$�����Q�-E�zW�l5n$�0��4WO�G&z��|��T�<��r��Xz�q�*���*i�В-L_O�B��pL����V����d��Gc]%��u���c��D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{����h�4i�)��a\�e1������)Xj�SL��t��v*�՟�_E�pI������1�Q,Z��I�6fD�������M���8%�t+2,>SU�P�r�����0�Μ�T>-+��$�|۷ �!����7^��\CT���GZ!&�]�����s���	)c��[D�b�1�,����O�r���Ҵ���;��B�yK~3,�RyV4 ��v�/�x��+CJ҆H/"U=4��"_wrhEc%A��� ��J A|�����|���W�w����N�]�吡�����C����'�M)�?Agχ[� G�ߑ�]�HF�K��ig|aj�'�)���p]������_�aF�q/Uolb�����N=���U�G�+��ZO�����v���5�y�	�󾈿Yp�)����[.-Zo|�;34���|��3��fx��D�Q��u$Vif���nO ])G}����P�0���Z�m����?�ܿ���Y�YHf�LB��sBH��|+%����s�-�IЫ���T���!�I�].��e�����O�S��70i�T{ �f�ch�j�v�Ta�Q����1W�>;+OXu�.n�Ne�����9ѵ���5�^�����P�C�7/�8V�R��k/�,YZU-,��z�7��7f.��ŤXj�=�#�2�6������'UO�K�4��c; 4��ژ@Z�0���ˬ�&�+�!Sw��C�꼵hEY� ^i~��_�����C8ܷ����9�˪�־�|5�m�������-A(�4\�Rq.z�?��h�{�����HMGHU�1�Z�q��}O�o�KƦ��H�&�i���D�$9W��c��7�	q��U��ns>E�
(9A�-tCc�2��`w�O?T�h1�
�R�i#ݞ������[�{C���?������`TX��f��^!�|�|s$����Y�¥@#k_�Ҕ2��u�\��I�N6ݳ&7}-p����s?�"E��2�t�I��#A`�}���M�s�͊��X���M��5+�:���/�4����!Wt�8�I"���"fp�:Kbŋ"O0��f���+_憔چޤֲ���A�8��Zz{�EI }��s��j�hH^Pw-{�ԪJy�X�o'OĈ�N�7'�]��c
w2�s��7�Ư�/x��kS�t��m�H��yϰ�V��j��q,U��dJO��P�;��%�T�I���D��h�+�/cD^��I�Ң����P	��[g\ћ{�{�g�9gt5\��"�"��_�����-�������Top�m-�0�&S|�nS3�%��9l�BK�Lۘ@w��n��H>�n;������.#�r�1��0�wP���"N� ~�O7��;2ԇ�SW���u$"[�1جU��y��.P���/�H�r12���� �^ˉя�}������j�k7��Z��)���L)&�.Q�ĆO�Q� A��8�&I����6I"��x��V�7�P R�2LR��33NH����gO��Q�^2��^��X՘���P� 6�W��@<��b��X�@�E4�V�|���^��Jb%Nf�������E&V(Wq8�Zr��$Wd<��#ֈ�Y��Dv����z_Y��Y*׏��xR-�頜�J�Vw-j�zB4�#�G	*��8�ު�M}��<鬘��{+���=z��O"���?�n�ʛ�2��c�l.�;c��fΰM���8FQ�j��>U�h6!Zؼ��$)��]	ӗj����>������8�:� ~-���j�J���_f+Y�t�@(1s�ŗ�U���/�a ��Fd�쉽�3�,���Z5鎟9����ɒ}�>��x�NN��؜���g�b����	U[J����(�N� i^筟��C|�9�Y����Ye]
L�)��&�����~���XP�!��R*�$Z)��6�� ���ݦ`�W1�a��u�08����3���K���{z� 0y���MQnSMS�&��wz�vF�����K�~����Qkj��`r"ub��y A+��x�R�n��q�Ov��+;�����>�'��pee���n�+
���1P�M=��% ��.��D���G�9���u��M���DNGʒ�]� �Ƅc�������Ƙs�ܡU�˒�)�x��YP/9�&t�)���`��|�G0F5�/���t���ۅ����v}�>�[�&��r}�:g��MI ����ρ�����p}����u��֪�F7���y�g:��W��v�N��6~n�b�A����gT�3$�d�Ŵ����<,N�;�u�眗�V|��'X�z��dDM ��4՗s�Ws�ݗم�m��Wf���1���tf3�-�`�w�z����[��ң�P5vxW�]�ch�)����l���ʝ��RK���8$L�`��Ҏ$}���!ּ�[�pއ�@4�?��hm�A�0�W	n|y:�t�wV<]�m��+.jI��h�����	�2����v��������끿w�@SP���yy�#���ݤI�P�p�p7ӫ?�m)�\5��E��w�����r�aYL��tI���<���jY��jU�J���`��5t��0�
���	>�[-w*$�=C��~[V��ܿ�˦v����2s��_�j���)DJp��σ0_�d��ނ�cn���*B8#�(��|�R��`�ۄr�޲n�F���.o� �8[*�ҹS_$ �
R��c�l�X�RD�_��sؼ��j�i��K9�>�_��3��n[۞���������ˏ��q7#��3�tW��O�6*���û'w�ze�@�]�U8�&h�O1Ѡ3��H1�r��.`��$����^#8��>W!*O���ͬ�5�:EdD>*:�9"�Q�g��z���(����m,�N���9H-Re^
��֩��c���r����үP����)7-�Q?���(��g�����N+�)�������7L��g�5
�a��E�4����r�������f�����)��3��'
����"ݕ<��Tpd|���Q��R�ϐɉU���h-�N��ؖ���t������^���-�>?T�p/���ܜ��Ck6�D���DW��X9�F�W+�^w]���I�撖6��}���M��P���Y�h-��`�u�dQ�n�!�R����&4�"��#��{hoLۧAnm+MD���	�/b��4��E^�W��?�����.0^`^dGUCt덮�螨�?E�����ȃh����Tw����q0�J�vy�4>x:�=�yryg��\K�^Γ�0ѳV|�x�WB��c�8.tqJ_�u 5���?���$ �5�*���$�#reY��rqђ���[�`�h�䬰*���In�d"J>F�a�-�:Cy媳�����Ay�{q�y�.�4`�QQ�������yʮ�����o>4�r���K�Ү���*�4>$�����g��l:b�O�U���(ePjV�ϕ���ǔ�a�}�]�K�����ٺ�X+�":}Mq>�}o���^LR���Snh�? ^���P�,�5F��3!�Y��'��f���gX��z1��!7�r���m�Ȥ 1�)��v`�#�x����e�2ެ*���r�~dx �I�/���&�"]8�v��t�$�Ͼ��7-��3܊����T�g."��^����� 3ew�R��Q����������6�#��ث���*���⟪@�ҧtI�m���ï�
�:d�J��j���f�TI#lA���j}����t3�#�g�$|\���3��N~6Ed�T�
:a����)�NYއ���s(&_
�孿���~�n4
p�BC��n��i
�&S��
%FX��Oy&�?b�G:��8Ad%����f��/��Q
�FD �lV��qֽ�X��\����)��RQ�ׄ������rLH����Zq����3��w{��zǝ9���YO���guԜ��k=��Omx���9�(�Y�Q��(mlNU-���P<��ay���Ql �Lw0�x�����Vd���d��K4೷V�04�tRS�ț�{	n����A娸��Y^�w�v�%'Lc	���l�2����1���eb1h���� �a먘�pؖR<5l�D�[^��!0H���F�D��(-yHJ�kY �����]��`�^!�P��%?�3z�(����@��KZ��b�{K�mgu� L���Ҏ�m�� ���HG
>f���
���U�^3_=��|�U���ROt�ע�4!2�T�"�_Y(~):u�TE'��!��ɢ'��_�D0�uR������X�B�	 L��4����('���b��M�"1+����t]��^�RM�>���f��D��]J0������:��/!ƥǌ� W����Wœ���=@o��c%M-�Iy�]�-}i��@Ŝ���Mrn���j����ۤ��'�HL*�+�'����!��O͂�+w8�@l�)���n`�:�V�p�ח-᤯M𙉵��J�?g�����1�]S[f��yzt+���R�v�mT
L�!�$���}��8�jkr�Y���X��*��,Mɡ\��f�bg'��GO��Q*U-�6c�;ľ�41�a�&q���k��|�C3�=GwD�6�9�B��JH8�c������L��NW��@�U'[���mǜ~n_T�#(.���1^o��$�mR�I2_tܐ�6FK䍸5SVb�n����o���A���p���sߓF��R�� �6�4��O��F��ʚ��I���\/�̓�ɯ-�ߐ�>�I��
ߎ�>̥[��DO�؏�� ���櫧�ٻ���1���.��pA�a�]�T�]��[H���!	&dƂyf���0�����|K������M%��.����]zbr����f$�YT����؀[%�����glv"֗ܕx�Ȼ�ɬ��#g	�`8x")��'����y\��j�LJ��o:}�^���3��g��l>>8\���J��Z���h��G}��"�Z�ٚ�b��i���{����s)b[DK9�e�O�,�<�!�Ȱ�3X�����W�1�44�,�2�^��^�6X���@���:e/��S+{۔�H�a���5����op�0���vl{dtO�}�8	p�'��7;�]u(Ef��D�D_Kߞ����X��zМ~�����ޥ]x$^7�o��vbXF&���u�_�v&�G�1��0Kߎ��OQ��ca�d���A���5<8#�ցV�^�D|�*��� �U.�;#�e!�Jj=$�c�D������r�m��n�&u�*�hc0ef+0�=�� ��7uЍ��"�}��9��v��*�dFuv�
�]�-����=2HJ5�Ѥ?�ۦ:_�mǳ���pN���qW��ݧ��C�v�E�~U08T=��8��"�y��*�O��K��B�T��[QQ�oG��6���eb¤��9^H�;��'��-�ݩ�q���#�-B���g2`9*���w&�]����'�_�ġ����=��J�*73֖Ⓔ�R��f��l�.2 sW�t�/VA|ZhcBrs�c�E��"y�˼ռ[w�U�i��I�ոR�?�}]����2��gD��ۚ���n��s1{ԃ@��B�Q�ؘ��p0|�Yҳ	D��刐�;Tc�����r�[,fڟZ(UR�T�����;���)�b�B{9����4f��,@�O�����$��7�}�8������Q{qv���3�e+�����O��9*��=����
�b*�-��G:Y��h�{�b{��҆҂�[�t=;��9�{5]�dO��X��c�����J�e��v�⬬MS�<�#���s�����|��	m�3��U=�?����i�v1:�Qj}�4KHf,�&�lk��xH��TM�!��p��F>���R��Kn��?��e����=l�J��B���K��$[ ��џ��#��"�`z_a�6$�9�[5eLF���i`��\0�*�+g���2sc*��bD�F�]V95Z� �*�Q�Eo�G�+hT�y��ń�K�HY�=!���E�^]a"�xP���X6tL�vW �"
*o~��X"}W+���#M&�B�o�y���ۓ�!!Y��T�P�4��*Pg��V���w�+�Sx����	�	�MqGj1�w�+Vd��]���'�u%w���=N�[>2�.��N�y>i�c�? <I����P��uѸ��.5�%ض�&�ZYa��^��r�h^ᰋ���(���[U��K�Zw��ɦn�(��4F��S�<�r��h�cT�0���hAkm��w+	_��� �;$k�%JwVaP!B����.��?�(�seOV���q����m��~ #�jrM��'�H��h�-��i��jǃ���fgH�#nQ��F�	e]N��>����5`	�Ʈ�_Lܥ�48+��	�&ĭ�N���Ŵ��d�Y�*]�^S/�y����ݵ�t�a�F��9�CFUy2,{H�Q܈��b�
��-�4Y���TrG-�B�Ʊ�G��JZ
Zv���P��3�o~�b�eD늫�xĴ�b��p���t����;������1�����Q�O��H|���}�4�B�G���I���`�8nB��}9Z���7��ا�`���P[��SZU�E��Gk0���#�y��0?Df��s��嵳⪦VP���5A�(Ц��M��|�mF�7Z�)=���+"��ے�P0� D�����5JF#'��.b5�<6�ѭ}#qҏ�	��x��4�KN��-J�n�~W/�{I���Tbژ�_r��h���9�ՠ���g���}o��a�ۍ�z:'���^C{�H ���LF�L~��iqB��6E4�Z�(
��D���7�g�ΪI��t{���L��J�;(��n��Py�)���S��JK���!4�C,�C�GZ+�7F����"b���ag�$����,������4�6��#*�@E��Ob�ð)��N�K���M�U�I\���԰����}J��tFD�#��|� �vƲ�n�Ux�S�I����{H o�M:"���M�"$��Z�`��1&|�����QkoC�5[���:icSA��3��9X߾���ұ������ah�_ y�/e�Df��sep=X�e?����:�2��a`�CH���+�U�g�՗΍�������7��#"��`�o�e�Iu���=���>�%�@�T'[�٪�3
=yqMB��iDbSs�P_��
hh�J�ȷ�z�w3�<�v�M�ԜR1.듅��Z��H_y�k�܂�v����*��/�~�O���;�q!�d~�L�3�U�Zf���ƙR�+�w�`��P�OL�.v�xK�'9+΢F����gwf�S"�-�N��
�j�����2t���u/~\���4�$̣���le����̽����`�{1oZ�zOMc�9� ���'�w㭺����dO�1a��kfƤ��0 ��o���Hm4�:��o�Dʓ����X��Ȍ�M�ܷ�I�x`�t��u[��2�Z7���5�� ��w��"���˧c�A�_cv/*�ڔ߬�}� Q'��
X=;�g��ԕ58���)g�f�1܎VȠ�C�}��?	�y�}�a���2��[����kL/[{d��Kɜ(�F3Z��Eo��͸�����j��m��
�֏9f�DTђE�zf:CBVI������l*].����B�D��l��d	�8�W:�{�ݞF�_� ��~���3�8�9[:�3nD8U�&>�x�k�ݔZ���6�7�g}G3z�����y��Z)X�-몳0�B�d�2EI�n�:�$f���D�Fpb�]3��i�$� �B�	uU��|��f�C�^��y���v-R�:'h'C����_]L���?��Ki�CY��(풕l�DA&%v�Wo�4�HӀXGi��G�r�pP��f�/���܇�U����x��u�q�kC�Mi�>\S��#qB$�t>��g�J�wv�T]m�4c��V����\4G�;�K_�Ƶ+6�ʶ���GO��-V���vs�fa��
��T=\V���+���n����я�Q�=�8���S}-����(1�2J� �0�i��BK��1kn�6���/b�&w��c�^nU��Ƴ���iܝ����l��C���6M�}�����@>U���m�+Ha�?��ڷN\�_���,W,����
P���pKR\t��]�?
b�'Cr���/���+��or��D'}Suj2����ț�	-L�������$3%(Ч�!9�T�K���q�b��<�02�v�\~4��q�����SR�*�-Ύ�5d�x^�/���Z�B��S#!��.����F�
x8�r�Y:�h�VV$vE`��A4��#eMsĠf k�ꃐ&��#��iK���9��4l_h�<ʃj�w��(��ѣad_�'bR�����m6V�����[��3a��X�P<����bS0򠱑F�r���)�M����&A��%��BO�m6
�2���lHff���¼u M��E���ӷM�K4�s�"#p�����/d�P��a�3�UP�Kj�U*k��zJ Q�|���E��>�����	��\�� d��w^.g����J����� Q���i	�Y��>��1�L�z�ۡC�j��/�q()Vt7N����b���į ��<�S-�闁 mm����cn0eT�3A��j�n�T2���DV��9����e��l*c�)+?d'��s��v���K���0�ӟËʧ�JA�m�d�R�`�!O <PA9u�&��E�KNP��&�ނ'��2�}��[�dg+��^�����F$��Z�}1{�6�^���[������"�˷��4��Ƽ~ҹV-?��i31�:��h����I�l�Ź���A/g�BM,zۃ������?a0��bJ ��Qz`v+ �\lTRJEJ�5���x�8p$�u>�ݐ�1�/ۺ�~�t�e��6���*�Ɠ�s�gg`��5�QF3���o

�2�nS�F� /�O�Kyuǵ�U#�� Y�1��l]�<�5��p��CŦsJ��I*�zT�%<��wz�+��O���9�&%"�����מ��Ô�-�R�wÌ�	.���Y8��x�ˠ�<r�K*t�92t�)e�Q���.��!�ID�\U�؅�+U���7�[���
yF�:f�亃N��GD���_ص�8B��Z~>G�b�M��yݟN%<���f���i��>����kd`NŎ�ሕ����n�K*��ޜX���.��~1ӹԣs[�p4�w��y�2'�u�����#n�(���
}�;@x��y�۞PG��g �B����x�e{��B3�����6�����3*��d֪�����1P@���`r��RWz>΍.��.4<���ck�|��7� B�k�	$Z.�eԧm�g��SlɵJ��[f ��C�P	پ��^��>�鵎`kR���L���]�yJ�z���f����89��j�8��O9&?"e��=<�S�T	�	YNE���WJ5��� ������Kf�W4Ċ�V��ʓTl8��~S$+I��P��G"����g#4W(��`��?	%���E#�&���0���D  X���wL�H(	TX�a=��	R��͐���OB�~!���-��ܦ��@�_i���i64W�cS_�Ԁ[�.�kJ�zj���H�fo���Q���"5��N��j�&��5�� ���`���1A��J)(��Ȣ5�&y���Ϸ�4T���%3�L���n�iq��1�뇿�i��k�*!KhO ����MG�y������@��_�M��]�`}T<XrVT	�Њ�l�(B"?�6z��DchƷw���,�ث�4��XAW�(�eK���A`FYر�Ր��S��#S7�B%	� 	��Ûȁ����5h.�W�4����7����-�7l���1��,ցz��]�K�K!=/�wV�F����y�+Q�N��;��i3�g�ܚ\"s��L6�}�)j��$�!�(F�7��Nj�B(
3a'�+�z����	ZBu�02�~��'��xgӁC��o|�4�<�{�^x��c_D������q�	��e�p�*Y�����������`X:���� S�T����3,^�^ �FL����@#�-�7L�u����݈�	X��è�i��Hu��zcՅ�Fև}�\�/wr�!��n@���4d�|��J�pI��Q^��5�!��|K�".�
(u��r>���*�$ɕ:�	M7�`��cx�Ġ,�V]#ϩ���a��#T��ݕfF���,J�({Y����<~��n�q�Y���Q��¨��A�I��F�w�嗠���l�"�I�T���-���Ɵ�F7l`�> ����������z���/Ǌ�ܫ|��&��\���c��dX�����[������ݵ�N{�4l��k���{8����+&b�S(8��O�� 8��Ξ���h��9�=�����a���:~���юp��>����D�-�O��+[Ҵ�n�\:L	�0.36��v���x���_��R����+�;ʌ��I�@��!�q,%��#=�	!�͐��ぴ\޽�O����m��������`Cc/|�.M|>I�՞�'�b�?D�){xƤ~�'�j	oY��¶��D��q��.�L�	�8ZП�G��k�����g(�7��L貅�q=�?��t&��ad�,ԧFj�,���yz:^��Ѳ@E�d�r���s�>\˜Ϗ��YM�t̴��j��{^&u8���8s|��3@�?�P�%5t�ٺ0D�g�0�sr��Q��֡�R�3ĭ��Vm��<x��#�@×�s��]�4�2S�̄Mb)��mu;�::�P���X�E�+z�;`�C^=������"#:Â�^:dU+J��H�苻���6*`�@��6�:G�-e�d5������_��p�@����7��䱉�Xf���Q}߃rF���b�JDw�'�~���zp�zY�G�~���O ���[��o�C�5�
����PTREP��p��_*ڸ��ȣ�y��g[)�:h`�U��:�v�X0��!��p�mDe\�u����G�ԉ��~# N^��N���D�R�ϲO=�ϼ�Ҹ9��8(�2Z9:���t=3�6_����Q�� �ԗڣ�����Cx�\��l۾�?	Ϸ9Rl�D/}6��堘8���'Ic�E�6��'wݳ��