��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��x���9eS� ]�_g�Xh3��1��63�A�1{Վ�eb��9��d8_��g�G�oWs$㩕�䫀�*Q���7е?-�@�Z��.޷�0�Ȭ�*
XL�1���-ec��D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E��,�׮ٴ�֘��w�{O�{C)\��z� �x=�ا�P�Bj0��d�	��-%!C��狎�{�]��� ���.w�C��ӿ^}E��V��{�0��GH�S��i��>	�R1H����l8i��<�������HIq��77}���/��� �5f2����_� Ыc���&��
V���_��:�D�X��rKJs#��i�k��B�y�����Ґ8�zC��V@D��j�Z�3?Z��m��9|b4�o��y�Z'�C��H���̍pL�BV��
Ö�=��/)��<S����Y	D��7���"DDB
|hK��@t�
K�l���;��ny@�%��uɁų�\�V-�_�*�v�wa����)�K����Cm�-k[�Z=��YTN!�J���+�y�0ܚ�4�ȹtŮ�ܣ`�3�����i�`�aʘ0�P;j偪�(sn��7�x�?QUY�*vg��X�:Mf��Ra6%%��2&��l��4�|.g���6W�e����% �|GKŻg��m�x	�t_A�t��v	�ԍB�Ǹ %�8��!��\�u�B��ˁR$vB����q07� ^ȣ-A��ϼ�o(�3�Pq�󲤎T7`�B'��`�狦����>�{<L��R[�G��ˠNfb&�ugo�g��.�� w����3R��k��]0$Aa�0S�M��\񨖄{6�R �B<��G4�SMŕ�շuo.m u�V�ZI��|U�׫썕�P�tf!#���riN�x>��\�����C�s�]�
M�h'�������p�|��Y�RҽO-Et��	�x*m�Vp1^�e�	�h['1+�}f��h��� 0Ǖ���Q�e;�/F���詣J"]��C�i��Wp��A]��'&w��]h>�A�"�UF���ѭ�f5�y��E��a��6 Hf0hɴ3.O�tJT�"P��*e��'�d��m��K����F�Q��ܰdk1^�Z�����1�W�kè�����#ǦR�0�Ŀ���9�J{`(emo���<��y�Q���}A8p֭x��཯��Ў�݀�q�&[�D�ܒ����K;I����h�jk���6 �ڦ���Jʳ {������)�I/W��k���Vy�=ӛ�M]����m\��8ϐ+�y��B�7ʡ��$֓l�i��n6�W�٭��m5vY`���x��QKf��nc+�
�Jnq2�#3	�o�̪��UwE�� ǯ��K�`�s�S��u��{��mY���Z��T�'�s6�<D�Ĳ�J9�S�A�c\��$�ڊ^��R�����A ����v4.��Y`�'�6?\�&j3d=25���'�e���,����j�xX�+Q���
��@��ť���BA1c��Jz� ����M諰8L�Y�r���mU���*Y��E��O��zw�NY
I]�W���|'q���Z�iK�W�gL�}h�7���`�*�
�K]�¨+��p�݆8��`A��ߍ�n/�f�um`y-��Y*�¦�׉�/���ړ�$��+h�}�xhY�$ ���A2Wgup
@�4���X`�����+S�Q��ʿm{�g�d3���8Q'tr�$IC���-�#w���.��hG��%�B�E��3wj�(G���_�ءpRח�tÖ��,�ǋ�@��76Ɯ�Vk �Ѐ�# Xd�Qg	g&{�5�����0��c� �*e�}c���dA�>��N�,7�d<w�|<w�1�l��X6gAj-FI��W�0�P��Lh�_Nƛ���� ����9n��]Q�?�$���N@ȣ�<��ub�ϫ8�˙J�-�`G��Tc���|U��u��_򼀆S�q`���6nmp��)��G���TYl)#���S\�Ƌ�E�(�͘1ǧ�z�Ag2}�eà4��:�}3������"G���4?�%��8��d�&MCQ�����Z������Yj�F_��;ۇGĜ����gNd|Ҳ1��������%����a u	�>�ʛ0�.O�l������҈p��U���
2�ކ*\�67N+8�M�a+��k�����Z>�![��'����|��
�p!��= 0Z�ki�����
L6R��e�;i��Ś����I�'���LE��1��z�9�4]�?��a��`�3[����R�e���Bd7t�3��J!�C9�D^�[@�5����訨2{h�%�鐨�!����<VV� cnGr���ON�~��E��sg���vz:6Q4� �?L�u�Fq���2�B�#�9p�NS$ nn�f�,	߰?62��i����ahA+nj����CNvFu+�i�����t:8V�����<=c.�x}��b2�5<�~w�c�.�t�OG2��oif�i�� oL�h7��@V��o���.�-�����D*1���+��"�6����_�Y���f=��8�S����p���+����1{�\ ���̇�XDҏBDt-an�P�J��v�R��%�.��1�MH�)���Mv�q�Sǵm��P�v�OL�,{,����8	��^�~�/� �c�#�|ω3�'\��#��@�T�>Ll��$L�.���W�A}���S�����:����a��F�)k
v��"J�g����3�[�uԟ����y͹W� �q��r��0^p�*�@�$��d��b��5��sz�npT$6�������;%��×6Ȣr�����/�*d��AF��[NK�Kl�����!²��l�DD�?_�C�����W�tA�@3~�і���i��%i�B�:@��9���1g��!�>�6 4�+Aj���%Z��`'�*B]���Ò���+W�����>H�ǘ������X����K�X�����T��nB��k<��Ji���hܻ��ٝ%�:�^��-eI__�[��q��gQX���a��O����[m��.;+���KR�؂i�P��ܼ��Awm���N�Ӊ�E��Nm?Ú4[`3WQ����3I��J���p?�*�^���;�mw	V�;��%'�S��2�yE�a,��Xw��T/�T�@��v6R�z�[��	j!H���?�%f|A��٠nl&�\�ǔ�$�>� �E������9����{v���7i�"��C���hD֠��b{�t.A�H�e6��Ġ��$��,����g��.����7k A����پ[�9�O�9+�FX��O_OvI152�r�ɱ9�-��92 �^�2u&���Z�5B�����s��-$zg]��L����c��au�/���eg(T�����Q���)���b>4�_&.��Cx�U�k� ����_rLh�0�DZ��|���)��D=J*&��)�y*-Q�U>I���-��'>x�����[�\��)^�Aě��3h�V�jv�Ve7e�֔��Re[���@`��?��zT��\�g������~5+��g���k>��:�X�n���߶���[d^�i��F�4��� �.��9�J{�ANH��qA�����n��n
��1(�s�iwE���9H�D �sp��AI�0a�qO��e���闍���*����� ؓg�����3`�*c>Z\˨8"oWi]{���KC8�Ը�h��.��2����²3��D9!`�N.5[l�eu^:��9(��{+'�0~�*g�ĕf~�(V�P��A����(4��:����lv�z���4�e��d`����ŧ<���>E<�s���cn�|N���N�2m*��<^J�G;k�w��0f�Zis ef6��G Զ�� �9�V=��a�[!��.�����K����ޛ/�*��a7�уîKv"> ű��S.�/�f�`f�%�ɳ��.k������m�)ㆶv��P�4�!�h\�����j�r�C�E_�@����wLآ���T�vt{$2J�P�R.g^l�p
6�%�l�+2��:�K"�_v��W�����O�{�G���m��\r�"��`�r^U�KE��r�q�{m�K�h��`�܈�d%��I��2����y��0��X3�v�a�2c��w��>�ӊ������vL
�� Z#����=��W�#�7M��W��³���!W8��7@VB��Y��D���$w~�"��Y��gG�@���?!m�
�E��Xi5�)�NX�F�
\[����U���Tﳣ�V�������ӵI9���񷮓i�<�V+Ş�l�
�i*yӷ8��"�