��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��x���9eS� ]�_g�Xh3��1��63�A�1{Վ�eb��9��d8_��g�G�oWs$㩕�䫀�*Q���7е?-�@�Z��.޷�0�Ȭ�*
XL�1���-ec��D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�9s��	��J�S��"�3�-��X��K���ȫGS$V�;�a.�DUzԖ�� ��>/XP�`��Q's�K"$�B��8��3�Ư����-��(cJ¸�qç��a�[T�e�W�[�G=�
\F��-���Xő	���GRA�[:KͿKB�S����������;@Eǭ��gŢF6�����w*ɓ�D�i�j'ۓ!��v殽	�3�^dujt�lg��$M�F��0B�A�u�w�$U7�!�N��������g���(p2S�{뽳�1󛉤־J��Z�D�%V���]k.���&�+e�d8�+N.L�Xme�?m�X��i�摉�ﱟ�9q�Oe7����m���%�T/�:�ޗp�
7�[���o�Z�rML���}�̸�d07�����\��E�� [���@��R �Ȯ�����8�&�є
Z`���ͯ84��U"E� ,��3����*r�0�ۀ�z^8�hb�08��O+�7�9I ͹0��FQ37Ğ�$�'���׌e��IڞG����>5�o�,�~
K�8��ؔ�Y"kƄY�.�ݏ@�O�1�/F���]y�}%�mYA7����Bƪ4�<I�'	���r}'5����"sN�A�ÿ�]��TH6��%��Ġ��� 釂�]O~a�޴�O��"a��9�7�*q�b����ݳr[Y����H�-�p=EW�2��2�1S��7�k�<"�����_�>[vm��%�
��25��W�d+5YJ�g~deA�w?$���[�:]��q�P�w��I���@��\ȇ�4����3H�ы�T��"��DDw��qQ�+<󽕇i��I�"��F��>u�s���^����E]�\�@}蓻WL¸ĸŦ{�;{��f�x4�tRi����w�����������\�{�n*�����i�|�)0	|bGƁ�W��`��GK#Y"WQ����N��Ŝ�l����?��~2uf>jLz��6Dr�o����3�őe�i���;�Z/B�Gb�C�w4��������<�W����[&��y`��3/m��H�͵��V���f`��H�oS 5:�X����o����G�3Է~w�i�j�\��pR��O]5��]`��£{�.%��dRK��}X(������ɺ�if �N?����3N��	a:b���,���Oj�YmT�GO3���]����s�ͱ󣃀����O=�us�уBA��)���h�M	ߓ>	���:�D��@�T-*('PO��#����|��Y�My�<��ݚ=�u0�����|٫F� ƻ��v��=�;/� ��e�+�Gȑ�,���Et��T���5Z���񧥵��!0>ho9�9L�%;�B�h���`�jqZ�N��{�/����˟�>)'KEɈ�fڦr�ƔO����J2� ��
E�d6�K=!yX4I?��h�qG���p[�A�{H�=��<MR,�Zr�өL79����妓��α/X�cu�`���N��Ր��j��_�Z2\������A�b@�K�R+��FS*L2SE��;��؁�i�j�[hZ+M%kɆ����=�������rO�4a�W ��7����;�y��m��E,n�v�\~Ms�!�5�Zu(�,�
ܑ�M��{�����n?,�ͼ~	���:�N������S~99��Vɩ	���F?zO��5��2)��0A���l�ī�lQ�N�X������vy���	k�;��q��=����Y��%�>�k�Wgyp"�{���Y5�m31HdD�s�8�(*�ܨ!%��G��
z�%7�Fc7�_�ŅUʣ�P��_z���vM^m�C�VԞ���z}���-�<KƋ��eZ�qah���{�F*>���x����1�.�#���Q�EG�}"��(�>ev�*L9$z�vT'y����U��_w���̈/睉�� �x=$��]��CH'g�l�r��7���������ʞ�7g�ou�e���.Os�3�v�OW^0f#����Ӛ��m��Fy��F�;o5�7�I����iC�_cR�C�A���9� ��1�<Wlxe�[q�#�+��ׇ���z& �j���b�fM~��ųSӞ'�	�<6�22��%ֲ�Y�fT����!rp�5^KBP1p����`o��3��-��P�R�@z֖B겚��9e�.f����#������΋��?��0;��*8P�<��n�a�} *�����8?` ���y���U�$甆=d�r�0��%�X����m$Yq�H�1����A<�_8BU�60�J�$�X�KO7��j��Z��zy?��)_=Uנ�6�����
m�[pBk�q�e%!��?z�G�*�J]�[rRW���.�_Cα�A���?WQ���}|��m���H!.�}�Bv��g�;��kQ'l���ᔓ�>85�A�����/2�W%eCx_�QL͂;0T��j���/#��U>����F��A�Qɮ�(:+�W�E���O��OY�@1�	v��_1�p�5��)�<c͕� ��b���,���*���&�v1��	K�+؆)#ӵ`�~�Qow�Kј��D��t���(yNL)����7	X��ŝ��x���\��R�g��\ۚ�H~�Ì	�][��>�ci�	�Y�����Z����D{��!���.��N�� �ӿ���ͦ�WiEWI�M
��b��{��?�y#��"*$x=��
 �c��Q^r��?��1:  �[��N�� �,I�4�8�R�e��w��Z0'����-�Loȅ�;�4愑m�[,���_�sWmg"G㭗�S�
c��"�C����u�ũT��r��9�3�l.<[g0e�%�c��Ό����k��#Uhj����\����@<,��%��C�d�z�S 囕g0�_�-R�j\��4/���W��p��t��c�]M���{���� ���("eax����z+4��f,N�N�N	p&����}�/��=��ȅ��BY&��"0gw)�.M?��>���N"Ņ�HU���F5���{V�c�H��f�#$yHy�Sk�n�>����z�4hC��	� &A�/N &���"ݺK-��Q���=�D�v��w���kU���;���z�b
�d�~�k�N��v���JX6����OV�E\��Mv?i�5E"KrsKI�Ɨ{�ȇ���r/�k.+@��;lR(֒rߕ��8�v�j{�bT{��i���NC�5fs�-w�M��vL��fg�H��8�N+n�,����,��X	Ռ�f�L�ʻC!���\�L����ve��Y�����c�T�G���� E�'k�_�Ыq���
A�9��Q:K�3����4���k�i[=�7C
���k����1�*�hT?�"����7y��-o���kS
�1,W��r��˃���W�I��Ԟ�L9�;������4^ػ#Kuz֞��&y���\�J����	څ2�p�K7����6����RQ>�7�X-x���Y��`z�s9�W���i�5���h�!�)�B���u��M=߉�M~ղ5+wط������@��,�C�_��U�M�E���M421"��36ހ7�獏$x�����?��sz��Ϟ�t8~ ���$�B�j��f�'�:��|)x��A�t�&��_2�^d;���i����_��>�3�.�CVE��ٯ=���#Ɵx�)ܭN��R�-1���e�:�%E9N�!�\�;��\a�b�d.	�b>��lSo�G�AV7��Ou���A�+�7g��V�L	;�����O
�uD�����$��?t4��i�tC?|�dx�����XE+8aؗ��Z7�����@�����7e���)��@-�<?�=x�B���E:�d�͓Q~�}�ɇ1m������}��3(v��g�<�<�3�K�����M30]t�1_��U���֋���VDZJ��M����� �F�yռqc8fH��Mo^X�,�ftJ��9�?<��f�<�!��5�����x�U�����Ds����b OS7Y.�	����=2g�ߕU�F����n7�^��`T!4�6��ϧ0<k��:��[Ji��c��I�r���!��E�@ւ�LF
�U�h>���ز�T�m�E�L�[�`9�٢�x�@צXQqpqR�CfX�l�h�d	�
+�����3�T���t�(�Ks�:�����#.Di�l�˨^�Vܼ���aa9�풡�r�p�;⇢�̫����읧j�V��1.�s�Ǒ��Rʎjʼ���/�h�yC�2�vvb�,�g5ż�)��>4�Ĺ�E�M������<,�_����(�R��E���C��7��|�l|��t�1��-�@y%F��eg�W]x����2�d��1~Ƙ���gm�7��7��-t�xȿ��#������"�3j9���s�r�*�Q���=�Ç��{�򭔝�*N5И�s�L��5-�	�f���Rɠ7���A��*�n�r]]��w�o=m��[�(ҷ|��̘��7�`
�55���I����v�O��0JW��\[a4��槩l���;��z5���`)<2�:{�<Р��%�;(�.L��3�\ŗ�iM/c��[���Zk �m�OL���g��e�2gA�'S
����z5��^Q�ĺ���5Đ� ��&߹,}u�|�%�W��=�jT%F4����{q����?���)